Spice deck to evaluate the static characteristics of CMOS, (W/L)p = 3(W/L)n

** Netlist description **

M1 out in vdd vdd pmos W = 1.125u L = 0.25u
M2 out in 0 0 nmos W = 0.375u L = 0.25u

cload out 0 10f
Vin in 0 2.5V
Vdd vdd 0 2.5V

** include library **

.LIB "tsmc_025um_model.mod.spice" cmos_models

** Static characteristics simulation commands **

.op 
.dc Vin 0 2.5 0.05

** Control/output commands

.control
run
setplot dc1
plot in out
.endc
.end
