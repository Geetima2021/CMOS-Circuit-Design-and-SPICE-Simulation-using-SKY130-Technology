Spice deck to plot the dynamic characteristics of cmos inverter circuit for wp/lp = 2wn/ln

*Model description
.param  temp = 27

*Netlist description
XM1 out in Vdd Vdd sky130_fd_pr__pfet_01v8 W = 0.84 L = 0.15
XM2 out in 0 0 sky130_fd_pr__nfet_01v8 W = 0.42 L = 0.15
cload out 0 10fF
Vin in 0 1.8V
Vdd Vdd 0 1.8V

*include model file
.lib "../../../sky130_fd_pr/models/sky130.lib.spice" ss

*simulation commands
.op
.dc Vin 0 1.8V 0.01

*interactive interpretor commandds
.control
run
display
setplot dc1
plot in out

.endc
.end
