Spice deck to find the dc characteristics of a CMOS inverter for wp/lp = 5wn/ln

*Model description
.param temp = 27

*Netlist description
XM1 out in Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2.1
XM2 out in 0 0 sky130_fd_pr__nfet_01v8 L=0.15 W=0.42
cload out 0 50fF
Vdd Vdd 0 1.8V
Vin in 0 1.8V

*include model file
.lib "../../../sky130_fd_pr/models/sky130.lib.spice" tt

*simulation commands
.op
.dc Vin 0 1.8V 0.01

*interactive interpretor commands
.control
run
display
setplot dc1
plot in out
.endc
.end
