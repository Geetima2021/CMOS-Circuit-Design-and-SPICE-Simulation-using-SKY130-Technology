Spice deck to plot the vtc characteristics of a cmos inverter circuit for wp/lp = wn/ln

** MODEL Description **
** NETLIST Description **

M1 out in vdd vdd pmos W = 0.375u L= 0.25u
M2 out in 0 0 nmos W = 0.375u L = 0.25u

cload out 0 10fF
Vin in 0 2.5V
Vdd vdd 0 2.5V

** SIMULATION COMMANDS **
.op
.dc Vin 0 2.5 0.05

** .include tsmc_025un_model.mod**
.lib "tsmc_025um_model.mod.spice" cmos_models

** interactive interpreter command
.control
run
setplot dc1
*display
plot in out 

.endc
.end
